library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 
 
package package2_2 is 
 
subtype my_logic is std_logic; 
 
end package2_2; 
